/*
 *  TOPPERS/HSP Kernel
 *      Toyohashi Open Platform for Embedded Real-Time Systems/
 *      High Reliable system Profile Kernel
 * 
 *  Copyright (C) 2008-2014 by Embedded and Real-Time Systems Laboratory
 *              Graduate School of Information Science, Nagoya Univ., JAPAN
 *  Copyright (C) 2012 by Ubiquitous Computing and Networking Laboratory
 *                Ritsumeikan Univ., JAPAN
 *
 *  �嵭����Ԥϡ��ʲ���(1)��(4)�ξ������������˸¤ꡤ�ܥ��եȥ���
 *  �����ܥ��եȥ���������Ѥ�����Τ�ޤࡥ�ʲ�Ʊ���ˤ���ѡ�ʣ������
 *  �ѡ������ۡʰʲ������ѤȸƤ֡ˤ��뤳�Ȥ�̵���ǵ������롥
 *  (1) �ܥ��եȥ������򥽡��������ɤη������Ѥ�����ˤϡ��嵭������
 *      ��ɽ�����������Ѿ�浪��Ӳ�����̵�ݾڵ��꤬�����Τޤޤη��ǥ���
 *      ����������˴ޤޤ�Ƥ��뤳�ȡ�
 *  (2) �ܥ��եȥ������򡤥饤�֥������ʤɡ�¾�Υ��եȥ�������ȯ�˻�
 *      �ѤǤ�����Ǻ����ۤ�����ˤϡ������ۤ�ȼ���ɥ�����ȡ�����
 *      �ԥޥ˥奢��ʤɡˤˡ��嵭�����ɽ�����������Ѿ�浪��Ӳ���
 *      ��̵�ݾڵ����Ǻܤ��뤳�ȡ�
 *  (3) �ܥ��եȥ������򡤵�����Ȥ߹���ʤɡ�¾�Υ��եȥ�������ȯ�˻�
 *      �ѤǤ��ʤ����Ǻ����ۤ�����ˤϡ����Τ����줫�ξ�����������
 *      �ȡ�
 *    (a) �����ۤ�ȼ���ɥ�����ȡ����Ѽԥޥ˥奢��ʤɡˤˡ��嵭����
 *        �ɽ�����������Ѿ�浪��Ӳ�����̵�ݾڵ����Ǻܤ��뤳�ȡ�
 *    (b) �����ۤη��֤��̤�������ˡ�ˤ�äơ�TOPPERS�ץ������Ȥ�
 *        ��𤹤뤳�ȡ�
 *  (4) �ܥ��եȥ����������Ѥˤ��ľ��Ū�ޤ��ϴ���Ū�������뤤���ʤ�»
 *      ������⡤�嵭����Ԥ����TOPPERS�ץ������Ȥ����դ��뤳�ȡ�
 *      �ޤ����ܥ��եȥ������Υ桼���ޤ��ϥ���ɥ桼������Τ����ʤ���
 *      ͳ�˴�Ť����ᤫ��⡤�嵭����Ԥ����TOPPERS�ץ������Ȥ�
 *      ���դ��뤳�ȡ�
 * 
 *  �ܥ��եȥ������ϡ�̵�ݾڤ��󶡤���Ƥ����ΤǤ��롥�嵭����Ԥ�
 *  ���TOPPERS�ץ������Ȥϡ��ܥ��եȥ������˴ؤ��ơ�����λ�����Ū
 *  ���Ф���Ŭ������ޤ�ơ������ʤ��ݾڤ�Ԥ�ʤ����ޤ����ܥ��եȥ���
 *  �������Ѥˤ��ľ��Ū�ޤ��ϴ���Ū�������������ʤ�»���˴ؤ��Ƥ⡤��
 *  ����Ǥ�����ʤ���
 * 
 *  @(#) $Id: kernel.cdl 945 2010-06-04 05:02:10Z ritsumei-takuya $
 */

/*
 *		TOPPERS/HRP2�����ͥ� ����ݡ��ͥ�ȵ��ҥե�����
 */

/*
 *  �����ͥ�Υ��󥯥롼�ɥե�����
 */
import_C("tecs_kernel.h");

/*
 *  ���������Τ�ƤӽФ�����Υ����˥���
 */
signature sTaskBody {
	void	main(void);
};

/*
 *  �������㳰�����롼�������Τ�ƤӽФ������˥���
 */
signature sTaskExceptionBody {
	void	main([in] TEXPTN pattern);
};

/*
 *  �����������뤿��Υ����˥���ʥ���������ƥ������ѡ�
 */
signature sTask {
	ER		activate(void);
	ER_UINT	cancelActivate(void);
	ER		terminate(void);
	ER		changePriority([in] PRI priority);
	ER		getPriority([out] PRI *p_priority);
	ER		refer([out] T_RTSK *pk_taskStatus);

	ER		wakeup(void);
	ER_UINT cancelWakeup(void);
	ER		releaseWait(void);
	ER		suspend(void);
	ER		resume(void);
	ER		raiseException([in] TEXPTN pattern);
    ER      referException([out] T_RTEX* pk_rtex);
    ER      startOverRunHandler([in] OVRTIM ovrtim);
    ER      stopOverRunHandler(void);
    ER      referOverRunHandler([out] T_ROVR *pk_rovr);
};

/*
 *  �����������뤿��Υ����˥�����󥿥�������ƥ������ѡ�
 */
[context("non-task")]
signature siTask {
	ER 		activate(void);
	ER		wakeup(void);
	ER		releaseWait(void);
	ER		raiseException([in] TEXPTN pattern);
    ER      disableWait(void);
    ER      enableWait(void);
    ER      startOverRunHandler([in] OVRTIM ovrtim);
    ER      stopOverRunHandler(void);
};

/*
 *  ������
 */
// =begin modified by ishikawa
[active, generate(HRP2TaskPlugin, "")]
celltype tTask {
	[inline]   entry	sTask	eTask;	/* ���������ʥ���������ƥ������ѡ�*/
	[inline]   entry	siTask	eiTask;	/* �����������󥿥�������ƥ������ѡ�*/
          	   call	sTaskBody	cBody;  /* ���������� */
    [optional] call	sTaskExceptionBody	cExceptionBody;
									/* �������㳰�����롼�������� */
	attr{
		ID				id = C_EXP("TSKID_$id$");
		/*
		 *  TA_NULL     0x00U   �ǥե������
		 * 	TA_ACT		0x01U	���������������˥�������ư����
		 */
		[omit] ATR		taskAttribute = C_EXP("TA_NULL");
		/*
		 * �������㳰�����롼����˻���Ǥ���°���Ϥʤ�����
		 * TA_NULL����ꤹ��
		 */
		[omit] ATR		exceptionAttribute = C_EXP("TA_NULL");
		[omit] PRI		priority;
        [omit] SIZE		stackSize = C_EXP("OMIT");
        [omit] SIZE		systemStackSize = C_EXP("OMIT");
        [omit] SIZE		userStackSize = C_EXP("OMIT");
        [omit] ACPTN    accessPattern[4] = { C_EXP("OMIT"), C_EXP("OMIT"), C_EXP("OMIT"), C_EXP("OMIT") };
	};

	FACTORY {
		/*
         * cfg�Ǥ�warning�����Τ���Υ�����
		 */
		write("tecsgen.cfg", "#include \"cb_type_only.h\"");
		write("cb_type_only.h", "#ifndef  TOPPERS_CB_TYPE_ONLY");
		write("cb_type_only.h", "#define  TOPPERS_CB_TYPE_ONLY");
		write("cb_type_only.h", "#endif   /*TOPPERS_CB_TYPE_ONLY*/");
		write("tecsgen.cfg", "#include \"$ct$_tecsgen.h\"");
		write("$ct$_factory.h", "#include \"kernel_cfg.h\"");
	};
};
// =end modified by ishikawa

/*
 *  ����������롼�������Τ�ƤӽФ�����Υ����˥���
 */
signature sInitializeRoutineBody {
	void	main(void);
};

/*
 *  ����������롼����
 */
[active, generate(HRP2HandlerPlugin, "INIT_ROUTINE")]
celltype tInitializeRoutine {
	call	sInitializeRoutineBody	cInitializeRoutine;
	
	attr {
		/*
		 * ����������롼����˻���Ǥ���°���Ϥʤ�����
		 * TA_NULL����ꤹ��
		 */
		[omit] ATR	attribute = C_EXP("TA_NULL");
	};

    /*
	factory {
		write("tecsgen.cfg",
			"ATT_INI({ %s, $cbp$, tInitializeRoutine_start });",
			attribute);
	};
    */
	FACTORY {
		write("tecsgen.cfg", "#include \"$ct$_tecsgen.h\"");
	};
};

/*
 *  ��λ�����롼�������Τ�ƤӽФ�����Υ����˥���
 */
signature sTerminateRoutineBody {
	void	main(void);
};

/*
 *  ��λ�����롼����
 */
[active, generate(HRP2HandlerPlugin, "TERM_ROUTINE")]
celltype tTerminateRoutine {
	call	sTerminateRoutineBody	cTerminateRoutine;

	attr {
		/*
		 * ��λ�����롼����˻���Ǥ���°���Ϥʤ�����
		 * TA_NULL����ꤹ��
		 */
		[omit] ATR	attribute = C_EXP("TA_NULL");
	};

    /*
	factory {
		write("tecsgen.cfg",
			"ATT_TER({ %s, $cbp$, tTerminateRoutine_start });",
			attribute);
	};
    */
	FACTORY {
		write("tecsgen.cfg", "#include \"$ct$_tecsgen.h\"");
	};
};


/*
 *  �ϥ�ɥ��ƤӽФ�����Υ����˥���
 */
[context("non-task")]
signature siHandlerBody {
	void   main(void);
};

/*
 *  ����ߥ����ӥ��롼����
 */
[active, generate(HRP2HandlerPlugin, "ISR")]
celltype tISR{
	call  siHandlerBody  ciBody;     /* ����ߥ����ӥ��롼��������*/

	attr {
		/*
		 * ����ߥ����ӥ��롼����˻���Ǥ���°���Ϥʤ�����
		 * TA_NULL����ꤹ��
		 */
		[omit] ATR   attribute = C_EXP( "TA_NULL" );
		[omit] INTNO interruptNumber;
		[omit] PRI   priority = 1;
	};

    /*
	factory{
		write("tecsgen.cfg", "ATT_ISR({ %s, $cbp$, %s, tISR_start, %s });",
			  attribute, interruptNumber, priority);
	};
    */
	FACTORY{
		write( "tecsgen.cfg", "#include \"$ct$_tecsgen.h\"" );
		write( "$ct$_factory.h", "#include \"kernel_cfg.h\"" );
	};

};


signature sConfigInterrupt{
	ER 		disable(void);
	ER 		enable(void);
};

/*
 *  ������׵�饤�� 
 */
[generate(HRP2HandlerPlugin, "CONFIG_INT")]
celltype tConfigInterrupt {
	[inline] entry sConfigInterrupt eConfigInterrupt;

	attr {
		INTNO interruptNumber;
		[omit] ATR   attribute =  C_EXP( "TA_NULL" );
		[omit] PRI   interruptPriority;
	};

    /*
	factory{
		write("tecsgen.cfg", "CFG_INT( %s,{ %s, %s});",
			  interruptNumber, attribute, interruptPriority);
	};
    */
};

/*
 *  ����ߥ����ӥ��롼����ȳ�����׵�饤���ʣ�祻�륿����
 */
[active]
composite tISRWithConfigInterrupt{
	entry sConfigInterrupt eConfigInterrupt;
	call  siHandlerBody  ciBody;     /* ����ߥ����ӥ��롼�������� */

	attr {
		/* ����ߥ����ӥ��롼���� */
		ATR   isrAttribute = C_EXP( "TA_NULL" );
		PRI   isrPriority = 1;
		INTNO interruptNumber;

		/* ������׵�饤�� */ 
		ATR   interruptAttribute =  C_EXP( "TA_NULL" );
		PRI   interruptPriority;
	};
	/* ����ߥ����ӥ��롼���� */
	cell tISR ISRMain{
		attribute = composite.isrAttribute;
		priority  = composite.isrPriority;
		interruptNumber = composite.interruptNumber;
		ciBody => composite.ciBody;
	};
	/* ������׵�饤�� */ 
	cell tConfigInterrupt ConfigInterrupt{
		interruptNumber = composite.interruptNumber;
		attribute = composite.interruptAttribute;
		interruptPriority = composite.interruptPriority;
	};
	composite.eConfigInterrupt => ConfigInterrupt.eConfigInterrupt;
};

/*
 *  �����ϥ�ɥ�����뤿��Υ����˥���ʥ���������ƥ������ѡ�
 */
signature sCyclic{
	ER 		start(void);
	ER 		stop(void);
	ER 		refer([out]T_RCYC *pk_cyclicHandlerStatus);
};

/*
 *  �����ϥ�ɥ�
 */
// =begin modified by ishikawa
// [active]
[active, generate(HRP2HandlerPlugin, "CYCLIC")]
celltype tCyclicHandler {
	[inline] entry sCyclic eCyclic; /* �����ϥ�ɥ�����ʥ���������ƥ������ѡ�*/
	call  siHandlerBody  ciBody;     /* �����ϥ�ɥ����� */

	attr {
		ID     id = C_EXP( "CYCHDLRID_$id$" );
		/*
		 *  TA_NULL     0x00U   �ǥե������
		 * 	TA_STA 		0x01U   �����ϥ�ɥ餬ư��Ƥ������
		 */
		[omit] ATR    attribute = C_EXP("TA_NULL");
		[omit] RELTIM cyclicTime;
		[omit] RELTIM cyclicPhase = 0;
        [omit] ACPTN  accessPattern[4] = { C_EXP("OMIT"), C_EXP("OMIT"), C_EXP("OMIT"), C_EXP("OMIT") };
	};

	FACTORY{
		write( "tecsgen.cfg", "#include \"$ct$_tecsgen.h\"" );
		write( "$ct$_factory.h", "#include \"kernel_cfg.h\"" );
	};
};
// =end modified by ishikawa

/*
 * �������򵯤��������ϥ�ɥ�ν���������
 */
celltype tCyclicTaskActivator{
	entry siHandlerBody eiBody;
	call  siTask        ciTask;
};

/*
 *  ����������
 */
[active]
composite tCyclicTask {
               entry sCyclic   eCyclic;/* �����ϥ�ɥ�����ʥ���������ƥ������ѡ�*/
               entry	sTask	eTask;	/* ���������ʥ���������ƥ������ѡ�*/
	           entry	siTask	eiTask;	/* �����������󥿥�������ƥ������ѡ�*/
	           call	sTaskBody	cBody;  /* ���������� */
    [optional] call	sTaskExceptionBody	cExceptionBody;
									/* �������㳰�����롼�������� */
	attr {
		/*
		 *  TA_NULL     0x00U   �ǥե������
		 * 	TA_STA 		0x01U   �����ϥ�ɥ餬ư��Ƥ������
		 */
		ATR    cyclicAttribute = C_EXP("TA_NULL");
		RELTIM cyclicTime;
		RELTIM cyclicPhase = 0;
		/*
		 * �������㳰�����롼����˻���Ǥ���°���Ϥʤ�����
		 * TA_NULL����ꤹ��
		 */
		ATR		exceptionAttribute = C_EXP("TA_NULL");
		PRI		priority;
		SIZE	stackSize;
	};
	cell tTask Task{
		/*
         * ��ư���˼�����������ư����������
         * ������������
		 * cyclicAttribute = C_EXP("TA_STA");�򵭽Ҥ���
		 */
		taskAttribute      = C_EXP("TA_NULL");
		exceptionAttribute = composite.exceptionAttribute;
		priority           = composite.priority;
		stackSize          = composite.stackSize;

		cBody => composite.cBody;
		cExceptionBody => composite.cExceptionBody;
	};
	cell tCyclicTaskActivator CyclicMain{
		ciTask = Task.eiTask;
	};
	cell tCyclicHandler CyclicHandler{
		ciBody = CyclicMain.eiBody;
		attribute = composite.cyclicAttribute;
		cyclicTime   = composite.cyclicTime;
		cyclicPhase  = composite.cyclicPhase;
	};
	composite.eTask   => Task.eTask;
	composite.eiTask  => Task.eiTask;
	composite.eCyclic => CyclicHandler.eCyclic;
};

/*
 *  ���顼��ϥ�ɥ�����뤿��Υ����˥���ʥ���������ƥ������ѡ�
 */
signature sAlarm{
	ER 		start([in] RELTIM alarmTime);
	ER 		stop(void);
    ER 		refer([out]T_RALM *pk_alarmStatus);
};

/*
 *  ���顼��ϥ�ɥ�����뤿��Υ����˥�����󥿥�������ƥ������ѡ�
 */
[context("non-task")]
signature siAlarm{
	ER 		start([in] RELTIM alarmTime);
	ER 		stop(void);
};

/*
 *  ���顼��ϥ�ɥ�
 */
// =begin modified by ishikawa
[active, generate(HRP2HandlerPlugin, "ALARM")]
celltype tAlarmHandler {
	[inline] entry sAlarm   eAlarm;     /* ���顼��ϥ�ɥ����ʥ���������ƥ������ѡ�*/
	[inline] entry siAlarm  eiAlarm;    /* ���顼��ϥ�ɥ���� ���󥿥�������ƥ������ѡ�*/
	call  siHandlerBody  ciBody;   /* ���顼��ϥ�ɥ����� */

	attr {
		ID     id = C_EXP( "ALMHDLRID_$id$" );
		/*
		 * ���顼��ϥ�ɥ�˻���Ǥ���°���Ϥʤ�����
		 * TA_NULL����ꤹ��
		 */
		[omit] ATR attribute = C_EXP("TA_NULL");
        [omit] ACPTN accessPattern[4] = { C_EXP("OMIT"), C_EXP("OMIT"), C_EXP("OMIT"), C_EXP("OMIT") };
	};

	FACTORY{
		write( "tecsgen.cfg", "#include \"$ct$_tecsgen.h\"" );
		write( "$ct$_factory.h", "#include \"kernel_cfg.h\"" );
	};
};
// =end modified by ishikawa

/*
 * ���ޥե��Υ����˥���ʥ���������ƥ������ѡ�
 */
signature sSemaphore{
	ER 		signal(void);
	ER 		wait(void);
	ER 		waitPolling(void);
	ER 		waitTimeout([in] TMO timeout);
	ER 		initialize(void);
	ER 		refer([out] T_RSEM *pk_semaphoreStatus);
};

/*
 *  ���ޥե��Υ����˥�����󥿥�������ƥ������ѡ�
 */
[context("non-task")]
signature siSemaphore {
	ER 		signal(void);
};
/*
 * ���ޥե��Υ��륿�������
 */
[generate(HRP2ObjectPlugin, "SEMAPHORE")]
celltype tSemaphore{

	[inline] entry  sSemaphore  eSemaphore;     /* ���ޥե����ʥ���������ƥ������ѡ�*/
	[inline] entry  siSemaphore eiSemaphore;    /* ���ޥե��ֵѡ��󥿥�������ƥ������ѡ�*/
	
	attr {
		ID      id = C_EXP( "SEMID_$id$" );
		[omit]  ATR attribute;
		[omit]  uint32_t count;
		[omit]  uint32_t max = 1;
		[omit]  ACPTN    accessPattern[4] = { C_EXP("OMIT"), C_EXP("OMIT"), C_EXP("OMIT"), C_EXP("OMIT") };
	};

	FACTORY{
		write( "$ct$_factory.h","#include \"kernel_cfg.h\"" );
	};
};

/*
 *  ���٥�ȥե饰�Υ����˥���ʥ���������ƥ������ѡ�
 */
signature sEventflag{
  	ER set([in] FLGPTN setPattern);
	ER clear([in] FLGPTN clearPattern);
  	ER wait([in] FLGPTN waitPattern, [in] MODE waitFlagMode, [out] FLGPTN *p_flagPattern);
	ER waitPolling([in] FLGPTN waitPattern, [in] MODE waitFlagMode, [out] FLGPTN *p_flagPattern);
	ER waitTimeout([in] FLGPTN waitPattern, [in] MODE waitFlagMode, [out] FLGPTN *p_flagPattern, [in] TMO timeout);
	ER initialize(void);
	ER refer([out]T_RFLG *pk_eventflagStatus);
};

/*
 *  ���٥�ȥե饰�Υ����˥�����󥿥�������ƥ������ѡ�
 */
[context("non-task")]
signature siEventflag {
	ER set([in] FLGPTN setPattern);
};
/*
 *  ���٥�ȥե饰
 */
[generate(HRP2ObjectPlugin, "EVENTFLAG")]
celltype tEventflag{
    
    [inline] entry  sEventflag  eEventflag;     /* ���٥�ȥե饰���ʥ���������ƥ������ѡ�*/
	[inline] entry  siEventflag eiEventflag;    /* ���٥�ȥե饰�����󥿥�������ƥ������ѡ�*/
	
	attr {
		ID      id = C_EXP( "FLGID_$id$" );
		/*
		 * TA_NULL �ǥե�����͡�FIFO�Ԥ���
         * TA_TPRI �Ԥ�����򥿥�����ͥ���ٽ�ˤ���
         * TA_WMUL ʣ���Υ��������ԤĤΤ����
         * TA_CLR  ���������Ԥ�������˥��٥�ȥե饰�򥯥ꥢ����
		 */
		[omit]  ATR attribute = C_EXP("TA_NULL");
		/*
		 * ���٥�ȥե饰�Υӥåȥѥ�����ν����
		 */
		[omit]  FLGPTN flagPattern;
        [omit]  ACPTN  accessPattern[4] = { C_EXP("OMIT"), C_EXP("OMIT"), C_EXP("OMIT"), C_EXP("OMIT") };
	};

	FACTORY{
		write( "$ct$_factory.h", "#include \"kernel_cfg.h\"" );
	};
};

/*
 *  �ǡ������塼�����뤿��Υ����˥���ʥ���������ƥ������ѡ�
 */
signature sDataqueue{
	ER 		send([in] intptr_t data);
	ER 		sendPolling([in] intptr_t data);
	ER 		sendTimeout([in] intptr_t data, [in]TMO timeout);
	ER 		sendForce([in] intptr_t data);
	ER 		receive([out] intptr_t *p_data);
	ER 		receivePolling([out] intptr_t *p_data);
	ER 		receiveTimeout([out] intptr_t *p_data, [in]TMO timeout);
	ER 		initialize(void);
	ER 		refer([out] T_RDTQ *pk_dataqueueStatus);
};

/*
 *  �ǡ������塼�����뤿��Υ����˥�����󥿥�������ƥ������ѡ�
 */
[context("non-task")]
signature siDataqueue {
	ER 		sendPolling([in] intptr_t data); 
	ER 		sendForce([in] intptr_t data);
};
/*
 *  �ǡ������塼
 */
[generate(HRP2ObjectPlugin, "DATAQUEUE")]
celltype tDataqueue {

	[inline] entry  sDataqueue  eDataqueue;     /* �ǡ������塼���ʥ���������ƥ������ѡ�*/
	[inline] entry  siDataqueue eiDataqueue;    /* �ǡ������塼�����󥿥�������ƥ������ѡ�*/
	
	attr {
		ID      id = C_EXP( "DTQID_$id$" );
		/*
		 * TA_NULL �ǥե�����͡�FIFO���
		 * TA_TPRI �����Ԥ�����򥿥�����ͥ���ٽ�ˤ���
		 */
		[omit] ATR     attribute = C_EXP( "TA_NULL" );
		[omit] uint_t  count = 1;
		[omit] void    *dtqmb = C_EXP( "NULL" );
		[omit] ACPTN   accessPattern[4] = { C_EXP("OMIT"), C_EXP("OMIT"), C_EXP("OMIT"), C_EXP("OMIT") };
	};

	FACTORY{
		write( "$ct$_factory.h","#include \"kernel_cfg.h\"" );
	};
};


/*
 *  ͥ���٥ǡ������塼�����뤿��Υ����˥���ʥ���������ƥ������ѡ�
 */
signature sPriorityDataqueue{
	ER 		send([in] intptr_t data, [in]PRI dataPriority);
	ER 		sendPolling([in] intptr_t data, [in]PRI dataPriority);
	ER 		sendTimeout([in] intptr_t data, [in]PRI dataPriority, [in]TMO timeout);
	ER 		receive([out] intptr_t *p_data, [out]PRI *p_dataPriority);
	ER 		receivePolling([out] intptr_t *p_data, [out]PRI *p_dataPriority);
 	ER 		receiveTimeout([out] intptr_t *p_data, [out]PRI *p_dataPriority,[in]TMO timeout);
	ER 		initialize(void);
	ER 		refer([out] T_RPDQ *pk_priorityDataqueueStatus);
};

/*
 *  ͥ���٥ǡ������塼�����뤿��Υ����˥�����󥿥�������ƥ������ѡ�
 */
[context("non-task")]
signature siPriorityDataqueue{
	ER 		sendPolling([in]intptr_t data, [in]PRI dataPriority);
};
/*
 *  ͥ���٥ǡ������塼
 */
[generate(HRP2ObjectPlugin, "PRIORITY_DATAQUEUE")]
celltype tPriorityDataqueue {
	[inline] entry  sPriorityDataqueue  ePriorityDataqueue;     /* ͥ���٥ǡ������塼���ʥ���������ƥ������ѡ�*/
	[inline] entry  siPriorityDataqueue eiPriorityDataqueue;    /* ͥ���٥ǡ������塼�����󥿥�������ƥ������ѡ�*/
	
	attr {
		ID      id = C_EXP( "PDTQID_$id$" );
		/*
		 * TA_NULL �ǥե�����͡�FIFO���
		 * TA_TPRI �����Ԥ�����򥿥�����ͥ���ٽ�ˤ���
		 */
		[omit] ATR     attribute = C_EXP( "TA_NULL" );
		[omit] uint_t  count = 1;       /* ͥ���٥ǡ������塼������ */
		[omit] PRI     maxDataPriority; /* ͥ���٥ǡ������塼�������Ǥ���ǡ���ͥ���٤κ����� */
		[omit] void    *pdqmb = C_EXP( "NULL" );/* ͥ���٥ǡ������塼�����ΰ����Ƭ���� */
		[omit] ACPTN   accessPattern[4] = { C_EXP("OMIT"), C_EXP("OMIT"), C_EXP("OMIT"), C_EXP("OMIT") };
	};

	FACTORY{
		write( "$ct$_factory.h","#include \"kernel_cfg.h\"" );
	};
};

/*
 *  ����Ĺ�������ס�������뤿��Υ����˥�����󥿥�������ƥ������ѡ�
 */
[deviate]
signature sFixedSizeMemoryPool{
	ER 		get([out] void **p_block);
	ER 		getPolling([out] void **p_block);
	ER 		getTimeout([out] void **p_block, [in] TMO timeout);
	ER 		release([in] const void *block);
	ER 		initialize(void);
	ER 		refer([out]T_RMPF *pk_memoryPoolFixedSizeStatus);
};

/*
 *  ����Ĺ����ס���
 */
[generate(HRP2ObjectPlugin, "FIXED_SIZE_MEMORYPOOL")]
celltype tFixedSizeMemoryPool{
	[inline] entry  sFixedSizeMemoryPool eFixedSizeMemoryPool; /* ����Ĺ����ס������ʥ���������ƥ������ѡ�*/
	
	attr {
		ID id = C_EXP( "MPFID_$id$" );
		/*
 		 * TA_NULL �ǥե�����͡�FIFO�Ԥ��� 
		 * TA_TPRI �Ԥ�����򥿥�����ͥ���ٽ�ˤ��� 
		 */
		[omit] ATR attribute = C_EXP("TA_NULL");
		[omit] uint32_t blockCount;
		[omit] uint32_t blockSize;
		[omit] MPF_T *mpf = C_EXP("NULL");
		/*����Ĺ����ס�������ΰ����Ƭ����*/
		[omit] void *mpfmb = C_EXP("NULL");
		[omit] ACPTN   accessPattern[4] = { C_EXP("OMIT"), C_EXP("OMIT"), C_EXP("OMIT"), C_EXP("OMIT") };
	};

	FACTORY{
		write( "$ct$_factory.h", "#include \"kernel_cfg.h\"" );
	};
};

[context("task")]
signature sKernel{

	ER		sleep(void);
	ER		sleepTimeout([in] TMO timeout);
	ER		delay([in] RELTIM delayTime);

	ER		exitTask(void);
	ER		getTaskId([out]ID *p_taskId);

	ER		rotateReadyQueue([in] PRI taskPriority);
	
	ER		getTime([out]SYSTIM *p_systemTime);
	ER		getMicroTime([out]SYSUTM *p_systemMicroTime);
	
	ER		lockCpu(void);
	ER		unlockCpu(void);
	ER		disableDispatch(void);
	ER		enableDispatch(void);
	ER      disableTaskException(void);
	ER      enableTaskException(void);
	ER      changeInterruptPriorityMask([in] PRI interruptPriority);
	ER      getInterruptPriorityMask([out] PRI *p_interruptPriority);

	ER		exitKernel(void);
	bool_t	senseContext(void);
	bool_t	senseLock(void);
	bool_t	senseDispatch(void);
	bool_t	senseDispatchPendingState(void);
	bool_t	senseKernel(void);
};

[context("non-task")]
signature siKernel {

	ER      getTaskId([out]ID *p_taskId);
	ER		rotateReadyQueue([in] PRI taskPriority);
	ER		getMicroTime([out]SYSUTM *p_systemMicroTime);
	
	ER      lockCpu(void);
	ER      unlockCpu(void);

	ER		exitKernel(void);
	bool_t	senseContext(void);
	bool_t	senseLock(void);
	bool_t	senseDispatch(void);
	bool_t	senseDispatchPendingState(void);
	bool_t	senseKernel(void);

	/* CPU�㳰�ϥ�ɥ���ǻ��Ѥ��� */
	bool_t	senseDispatchPendingStateCPU([in] const void * p_exceptionInfomation);
	bool_t	senseTaskExceptionPendingStateCPU([in] const void * p_exceptionInfomation);
};

//[singleton, generate(HRP2KernelObjectPlugin, "")]
[singleton, generate(HRP2ObjectPlugin, "KERNEL")]
celltype tKernel{

	[inline] entry sKernel  eKernel;
	[inline] entry siKernel eiKernel;
	attr {
        [omit] ACPTN   accessPattern[4] = { C_EXP("OMIT"), C_EXP("OMIT"), C_EXP("OMIT"), C_EXP("OMIT") };
    };
};

// =begin added by ishikawa
signature sMessageBuffer{
    ER send([in, size_is(size)] const uint8_t* message, [in] uint32_t size);
    ER sendPolling([in, size_is(size)] const uint8_t *message, 
                   [in] uint32_t size);
    ER sendTimeout([in, size_is(size)] const uint8_t *message, 
                   [in] uint32_t size, [in] TMO timeout);
    ER_UINT receive([out] uint8_t *message);
    ER_UINT receivePolling([out] uint8_t *message);
    ER_UINT receiveTimeout([out] uint8_t *message, [in] TMO timeout);
    void initialize(void);
    ER refer([out] T_RMBF *packet);
};

[generate(HRP2ObjectPlugin, "MESSAGE_BUFFER")]
celltype tMessageBuffer{
	[inline] entry sMessageBuffer eMessageBuffer;
  
	attr {
		ID      id = C_EXP( "MBFID_$id$" );
        /*
         * �����Ԥ����塼����³���
         * TA_NULL: FIFO
         * TA_TPRI: ͥ���ٽ�
         */
        [omit]  ATR attribute = C_EXP("TA_NULL");
		[omit]  uint32_t maxSize;
		[omit]  uint32_t bufferSize;
		[omit]  void *mbfmb = C_EXP("NULL");
		[omit]  ACPTN    accessPattern[4] = { C_EXP("OMIT"), C_EXP("OMIT"), C_EXP("OMIT"), C_EXP("OMIT") };
	};

	FACTORY{
		write( "$ct$_factory.h","#include \"kernel_cfg.h\"" );
	};
};
// =end added by ishikawa
