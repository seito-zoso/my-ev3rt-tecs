/*
 *  tEV3Sample.cdl
 *
 *  VM$B$N8D?t$K1~$8$F(BCDL$B%U%!%$%k$rA*Br$9$k(B
 *  (VM$B$r#2$D;H$&>l9g!$(BVM2.cdl$B$r%$%s%]!<%H$9$k!K(B
 *
 */
const int32_t MRUBY_VM_STACK_SIZE = 81920;

//import("VM1_bigtire.cdl");
import("VM2_bigtire.cdl");
