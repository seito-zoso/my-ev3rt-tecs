/*
 *  Copyright (C) 2013 by Embedded and Real-Time Systems Laboratory
 *              Graduate School of Information Science, Nagoya Univ., JAPAN
 *  Copyright (C) 2013 by Ubiquitous Computing and Networking Laboratory
 *              Ritsumeikan Univ., JAPAN
 *  Copyright (C) 2014 by Osaka Univ., JAPAN
 *
 *  上記著作権者は，以下の(1)〜(4)の条件を満たす場合に限り，本ソフトウェ
 *  ア（本ソフトウェアを改変したものを含む．以下同じ）を使用・複製・改
 *  変・再配布（以下，利用と呼ぶ）することを無償で許諾する．
 *  (1) 本ソフトウェアをソースコードの形で利用する場合には，上記の著作
 *      権表示，この利用条件および下記の無保証規定が，そのままの形でソー
 *      スコード中に含まれていること．
 *  (2) 本ソフトウェアを，ライブラリ形式など，他のソフトウェア開発に使
 *      用できる形で再配布する場合には，再配布に伴うドキュメント（利用
 *      者マニュアルなど）に，上記の著作権表示，この利用条件および下記
 *      の無保証規定を掲載すること．
 *  (3) 本ソフトウェアを，機器に組み込むなど，他のソフトウェア開発に使
 *      用できない形で再配布する場合には，次のいずれかの条件を満たすこ
 *      と．
 *    (a) 再配布に伴うドキュメント（利用者マニュアルなど）に，上記の著
 *        作権表示，この利用条件および下記の無保証規定を掲載すること．
 *    (b) 再配布の形態を，別に定める方法によって，TOPPERSプロジェクトに
 *        報告すること．
 *  (4) 本ソフトウェアの利用により直接的または間接的に生じるいかなる損
 *      害からも，上記著作権者およびTOPPERSプロジェクトを免責すること．
 *      また，本ソフトウェアのユーザまたはエンドユーザからのいかなる理
 *      由に基づく請求からも，上記著作権者およびTOPPERSプロジェクトを
 *      免責すること．
 *
 *  本ソフトウェアは，無保証で提供されているものである．上記著作権者お
 *  よびTOPPERSプロジェクトは，本ソフトウェアに関して，特定の使用目的
 *  に対する適合性も含めて，いかなる保証も行わない．また，本ソフトウェ
 *  アの利用により直接的または間接的に生じたいかなる損害に関しても，そ
 *  の責任を負わない．
 *
 *  @(#) $Id: tButton.cdl 5 2014-10-29 19:06:11Z hopf-takuya $
 */
import_C("ff.h");

signature sFatFile {
 /* ファイルアクセス */ /* void -> TCHAR に変更 */
  // FRESULT fopen ([in,string] const TCHAR* path_new, [in] BYTE mode); /* Open or create a file */
  FRESULT fopen ([in,string] const TCHAR* path, [in,string] const TCHAR* mode); /* Open or create a file */
  FRESULT fclose (void);         /* Close an open file object */
  FRESULT fread ([out,size_is(btr)] TCHAR* buffer, [in] UINT btr);  /* Read data from a file */
  FRESULT fwrite ([in,size_is(btw)] const TCHAR* buffer, [in] UINT btw, [out] UINT* bw);   /* Write data to a file */
  // FRESULT forward ([in] const FIL* fp, [in] UINT(*func)(const BYTE*,UINT), [in] UINT btf, [out] UINT* bf); /* Forward data to the stream */
  // FRESULT lseek ([in] const FIL* fp, [in] DWORD ofs); /* Move file pointer of a file object */
  // FRESULT truncate ([in] const FIL* fp);                   /* Truncate file */
  // FRESULT sync ([in] const FIL* fp);                     /* Flush cached data of a writing file */
  // int putc ([in] TCHAR chr, [in] const FIL* fp);                    /* Put a character to the file */
  // int puts ([in,string] const TCHAR* str, [in] const FIL* cp);               /* Put a string to the file */
  // // int printf ([in] FIL* fp, [in] const TCHAR* str, ...);            /* Put a formatted string to the file */
  // // TCHAR* gets (TCHAR* buff, int len, FIL* fp);
/* ファイル/ディレクトリ管理 */
  // FRESULT mkdir ([in,string] const TCHAR* path);                /* Create a sub directory */
  // FRESULT unlink ([in,string] const TCHAR* path);               /* Delete an existing file or directory */
  // FRESULT rename ([in,string] const TCHAR* path_old, [in,string] const TCHAR* path_new);  /* Rename/Move a file or directory */
  // FRESULT stat ([in,string] const TCHAR* path, [out] FILINFO* fno);         /* Get file status */
  // FRESULT chmod ([in,string] const TCHAR* path, [in] BYTE value, [in] BYTE mask);     /* Change attribute of the file/dir */
  // FRESULT utime ([in,string] const TCHAR* path, [in] const FILINFO* fno);      /* Change times-tamp of the file/dir */
  // FRESULT chdir ([in,string] const TCHAR* path);                /* Change current directory */
  // FRESULT chdrive ([in,string] const TCHAR* path);                /* Change current drive */
  // FRESULT getcwd ([out,string] TCHAR* buff, [in] UINT len);             /* Get current directory */
/* ボリューム管理 */
  // FRESULT getlabel ([in,string] const TCHAR* path, [out,string] TCHAR* label, [out] DWORD* vsn); /* Get volume label */
  // FRESULT setlabel ([in,string] const TCHAR* label);              /* Set volume label */
  // FRESULT mkfs ([in,string] const TCHAR* path, [in] BYTE sfd, [in] UINT au);        /* Create a file system on the volume */
  // // FRESULT fdisk ([in] BYTE pdrv, [in] const DWORD szt[], [in] void* work);     /* Divide a physical drive into some partitions */
};


celltype tFatFile {
  entry sFatFile eFatFile;
  var {
    FIL fs; /* ファイルポインタ */
    // UINT bw; /* write 書き込まれたバイト数を格納する */
    UINT br; /* read 読みだされたバイト数を格納する */
    TCHAR read_buff[100]; /* read 読み出したデータを格納するバッファ */
  };
};
