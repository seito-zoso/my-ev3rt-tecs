/*
 *  tReceive.cdl
 *
 *
 */
import("tFatFile.cdl");
import(<mruby.cdl>);
// import(<sMruby.cdl>);
// import(<tTLSFMalloc.cdl>);
// import("tFatFile.cdl");

signature sReceive {
  void receive ([in,string] const char_t* path);
};

/*** tReceive ***/
celltype tReceive {
  entry sReceive eReceive;
  call sFatFile cFatFile;
  /* MrubyBridgePlugin の生成する VM_TECSInitializeer.eInitialize へ結合する */
  [optional]  call nMruby::sInitializeBridge cInit;
  attr {
    [omit]char_t *mrubyLib;
    //[omit]char_t *mrubyApp;
    uint8_t *irepLib     = C_EXP("&$cell_global$_irep");
    uint32_t irepAppSize = 131072;
    // FLGPTN setptn;
  };
  var {
      mrb_state *mrb;
      mrbc_context *context;
      [size_is(irepAppSize)] uint8_t *irepApp; // __attribute__((nocommon));
      [size_is(irepAppSize)] uint16_t *bw;
      FIL fs;
  };

    factory{
      write("Makefile.tecsgen", "POST_TECSGEN_TARGET := $(POST_TECSGEN_TARGET) $cell_global$_mrb.c");
      write("Makefile.tecsgen", "$cell_global$_mrb.c : %s tecs.timestamp Makefile", mrubyLib);
      write("Makefile.tecsgen", "	$(MRBC) -B$cell_global$_irep -o$cell_global$_mrb.c %s", mrubyLib);
      write("Makefile.tecsgen", "TECS_COBJS := $(TECS_COBJS) $cell_global$_mrb.o");
      write("Makefile.tecsgen", "MRB_C := $(MRB_C) $cell_global$_mrb.c");
      write("$ct_global$_factory.h","extern const char_t *$cell_global$_irep;");
    };
};
