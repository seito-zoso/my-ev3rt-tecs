/*
 *   RiteVM$B%9%1%8%e!<%i$N%;%k%?%$%W5-=R(B
 */
celltype tRiteVMSchedulerMain{
    require tKernel.eiKernel;
    entry siHandlerBody eiBody;
    
    attr {
        PRI priority;
	};
};

[active]
composite tRiteVMScheduler {
    attr {
		/*
		 *  TA_NULL     0x00U   $B%G%U%)%k%HCM(B
		 * 	TA_STA 		0x01U   $B<~4|%O%s%I%i$,F0:n$7$F$$$k>uBV(B
		 */
        ATR    cyclicAttribute = C_EXP("TA_NULL");
        RELTIM cyclicTime = 1;  /* $B<~4|;~4V(B */
        RELTIM cyclicPhase = 1;
    };

    cell tRiteVMSchedulerMain RiteVMSchedulerMain{
        priority = C_EXP("RITEVM_PRIORITY");
    };
    cell tCyclicHandler CyclicHandler{
        ciBody = RiteVMSchedulerMain.eiBody;
        attribute = composite.cyclicAttribute;
        cyclicTime = composite.cyclicTime;
        cyclicPhase = composite.cyclicPhase;
    };
};
